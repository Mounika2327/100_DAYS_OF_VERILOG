module xor_gate (
    input wire a,  // Input a
    input wire b,  // Input b
    output wire y  // Output y
);

    // XOR operation
    assign y = a ^ b;

endmodule
