module not_gate (
    input wire a,  // Input a
    output wire y  // Output y
);

    // NOT operation
    assign y = ~a;

endmodule
